module GRReg(
  input         clock,
  input         reset,
  output [63:0] io_ALU_GRReg_IO_rj,
  output [63:0] io_ALU_GRReg_IO_rk,
  output [63:0] io_ALU_GRReg_IO_rd_in,
  input  [63:0] io_ALU_GRReg_IO_rd,
  input  [31:0] io_rj_addr,
  input  [31:0] io_rk_addr,
  input  [31:0] io_rd_addr
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [63:0] _RAND_12;
  reg [63:0] _RAND_13;
  reg [63:0] _RAND_14;
  reg [63:0] _RAND_15;
  reg [63:0] _RAND_16;
  reg [63:0] _RAND_17;
  reg [63:0] _RAND_18;
  reg [63:0] _RAND_19;
  reg [63:0] _RAND_20;
  reg [63:0] _RAND_21;
  reg [63:0] _RAND_22;
  reg [63:0] _RAND_23;
  reg [63:0] _RAND_24;
  reg [63:0] _RAND_25;
  reg [63:0] _RAND_26;
  reg [63:0] _RAND_27;
  reg [63:0] _RAND_28;
  reg [63:0] _RAND_29;
  reg [63:0] _RAND_30;
  reg [63:0] _RAND_31;
  reg [63:0] _RAND_32;
  reg [63:0] _RAND_33;
  reg [63:0] _RAND_34;
  reg [63:0] _RAND_35;
  reg [63:0] _RAND_36;
  reg [63:0] _RAND_37;
  reg [63:0] _RAND_38;
  reg [63:0] _RAND_39;
  reg [63:0] _RAND_40;
  reg [63:0] _RAND_41;
  reg [63:0] _RAND_42;
  reg [63:0] _RAND_43;
  reg [63:0] _RAND_44;
  reg [63:0] _RAND_45;
  reg [63:0] _RAND_46;
  reg [63:0] _RAND_47;
  reg [63:0] _RAND_48;
  reg [63:0] _RAND_49;
  reg [63:0] _RAND_50;
  reg [63:0] _RAND_51;
  reg [63:0] _RAND_52;
  reg [63:0] _RAND_53;
  reg [63:0] _RAND_54;
  reg [63:0] _RAND_55;
  reg [63:0] _RAND_56;
  reg [63:0] _RAND_57;
  reg [63:0] _RAND_58;
  reg [63:0] _RAND_59;
  reg [63:0] _RAND_60;
  reg [63:0] _RAND_61;
  reg [63:0] _RAND_62;
  reg [63:0] _RAND_63;
`endif // RANDOMIZE_REG_INIT
  reg [63:0] GRReg_0; // @[GRReg.scala 22:24]
  reg [63:0] GRReg_1; // @[GRReg.scala 22:24]
  reg [63:0] GRReg_2; // @[GRReg.scala 22:24]
  reg [63:0] GRReg_3; // @[GRReg.scala 22:24]
  reg [63:0] GRReg_4; // @[GRReg.scala 22:24]
  reg [63:0] GRReg_5; // @[GRReg.scala 22:24]
  reg [63:0] GRReg_6; // @[GRReg.scala 22:24]
  reg [63:0] GRReg_7; // @[GRReg.scala 22:24]
  reg [63:0] GRReg_8; // @[GRReg.scala 22:24]
  reg [63:0] GRReg_9; // @[GRReg.scala 22:24]
  reg [63:0] GRReg_10; // @[GRReg.scala 22:24]
  reg [63:0] GRReg_11; // @[GRReg.scala 22:24]
  reg [63:0] GRReg_12; // @[GRReg.scala 22:24]
  reg [63:0] GRReg_13; // @[GRReg.scala 22:24]
  reg [63:0] GRReg_14; // @[GRReg.scala 22:24]
  reg [63:0] GRReg_15; // @[GRReg.scala 22:24]
  reg [63:0] GRReg_16; // @[GRReg.scala 22:24]
  reg [63:0] GRReg_17; // @[GRReg.scala 22:24]
  reg [63:0] GRReg_18; // @[GRReg.scala 22:24]
  reg [63:0] GRReg_19; // @[GRReg.scala 22:24]
  reg [63:0] GRReg_20; // @[GRReg.scala 22:24]
  reg [63:0] GRReg_21; // @[GRReg.scala 22:24]
  reg [63:0] GRReg_22; // @[GRReg.scala 22:24]
  reg [63:0] GRReg_23; // @[GRReg.scala 22:24]
  reg [63:0] GRReg_24; // @[GRReg.scala 22:24]
  reg [63:0] GRReg_25; // @[GRReg.scala 22:24]
  reg [63:0] GRReg_26; // @[GRReg.scala 22:24]
  reg [63:0] GRReg_27; // @[GRReg.scala 22:24]
  reg [63:0] GRReg_28; // @[GRReg.scala 22:24]
  reg [63:0] GRReg_29; // @[GRReg.scala 22:24]
  reg [63:0] GRReg_30; // @[GRReg.scala 22:24]
  reg [63:0] GRReg_31; // @[GRReg.scala 22:24]
  reg [63:0] GRReg_32; // @[GRReg.scala 22:24]
  reg [63:0] GRReg_33; // @[GRReg.scala 22:24]
  reg [63:0] GRReg_34; // @[GRReg.scala 22:24]
  reg [63:0] GRReg_35; // @[GRReg.scala 22:24]
  reg [63:0] GRReg_36; // @[GRReg.scala 22:24]
  reg [63:0] GRReg_37; // @[GRReg.scala 22:24]
  reg [63:0] GRReg_38; // @[GRReg.scala 22:24]
  reg [63:0] GRReg_39; // @[GRReg.scala 22:24]
  reg [63:0] GRReg_40; // @[GRReg.scala 22:24]
  reg [63:0] GRReg_41; // @[GRReg.scala 22:24]
  reg [63:0] GRReg_42; // @[GRReg.scala 22:24]
  reg [63:0] GRReg_43; // @[GRReg.scala 22:24]
  reg [63:0] GRReg_44; // @[GRReg.scala 22:24]
  reg [63:0] GRReg_45; // @[GRReg.scala 22:24]
  reg [63:0] GRReg_46; // @[GRReg.scala 22:24]
  reg [63:0] GRReg_47; // @[GRReg.scala 22:24]
  reg [63:0] GRReg_48; // @[GRReg.scala 22:24]
  reg [63:0] GRReg_49; // @[GRReg.scala 22:24]
  reg [63:0] GRReg_50; // @[GRReg.scala 22:24]
  reg [63:0] GRReg_51; // @[GRReg.scala 22:24]
  reg [63:0] GRReg_52; // @[GRReg.scala 22:24]
  reg [63:0] GRReg_53; // @[GRReg.scala 22:24]
  reg [63:0] GRReg_54; // @[GRReg.scala 22:24]
  reg [63:0] GRReg_55; // @[GRReg.scala 22:24]
  reg [63:0] GRReg_56; // @[GRReg.scala 22:24]
  reg [63:0] GRReg_57; // @[GRReg.scala 22:24]
  reg [63:0] GRReg_58; // @[GRReg.scala 22:24]
  reg [63:0] GRReg_59; // @[GRReg.scala 22:24]
  reg [63:0] GRReg_60; // @[GRReg.scala 22:24]
  reg [63:0] GRReg_61; // @[GRReg.scala 22:24]
  reg [63:0] GRReg_62; // @[GRReg.scala 22:24]
  reg [63:0] GRReg_63; // @[GRReg.scala 22:24]
  wire [63:0] _GEN_1 = 6'h1 == io_rj_addr[5:0] ? GRReg_1 : GRReg_0; // @[GRReg.scala 24:{24,24}]
  wire [63:0] _GEN_2 = 6'h2 == io_rj_addr[5:0] ? GRReg_2 : _GEN_1; // @[GRReg.scala 24:{24,24}]
  wire [63:0] _GEN_3 = 6'h3 == io_rj_addr[5:0] ? GRReg_3 : _GEN_2; // @[GRReg.scala 24:{24,24}]
  wire [63:0] _GEN_4 = 6'h4 == io_rj_addr[5:0] ? GRReg_4 : _GEN_3; // @[GRReg.scala 24:{24,24}]
  wire [63:0] _GEN_5 = 6'h5 == io_rj_addr[5:0] ? GRReg_5 : _GEN_4; // @[GRReg.scala 24:{24,24}]
  wire [63:0] _GEN_6 = 6'h6 == io_rj_addr[5:0] ? GRReg_6 : _GEN_5; // @[GRReg.scala 24:{24,24}]
  wire [63:0] _GEN_7 = 6'h7 == io_rj_addr[5:0] ? GRReg_7 : _GEN_6; // @[GRReg.scala 24:{24,24}]
  wire [63:0] _GEN_8 = 6'h8 == io_rj_addr[5:0] ? GRReg_8 : _GEN_7; // @[GRReg.scala 24:{24,24}]
  wire [63:0] _GEN_9 = 6'h9 == io_rj_addr[5:0] ? GRReg_9 : _GEN_8; // @[GRReg.scala 24:{24,24}]
  wire [63:0] _GEN_10 = 6'ha == io_rj_addr[5:0] ? GRReg_10 : _GEN_9; // @[GRReg.scala 24:{24,24}]
  wire [63:0] _GEN_11 = 6'hb == io_rj_addr[5:0] ? GRReg_11 : _GEN_10; // @[GRReg.scala 24:{24,24}]
  wire [63:0] _GEN_12 = 6'hc == io_rj_addr[5:0] ? GRReg_12 : _GEN_11; // @[GRReg.scala 24:{24,24}]
  wire [63:0] _GEN_13 = 6'hd == io_rj_addr[5:0] ? GRReg_13 : _GEN_12; // @[GRReg.scala 24:{24,24}]
  wire [63:0] _GEN_14 = 6'he == io_rj_addr[5:0] ? GRReg_14 : _GEN_13; // @[GRReg.scala 24:{24,24}]
  wire [63:0] _GEN_15 = 6'hf == io_rj_addr[5:0] ? GRReg_15 : _GEN_14; // @[GRReg.scala 24:{24,24}]
  wire [63:0] _GEN_16 = 6'h10 == io_rj_addr[5:0] ? GRReg_16 : _GEN_15; // @[GRReg.scala 24:{24,24}]
  wire [63:0] _GEN_17 = 6'h11 == io_rj_addr[5:0] ? GRReg_17 : _GEN_16; // @[GRReg.scala 24:{24,24}]
  wire [63:0] _GEN_18 = 6'h12 == io_rj_addr[5:0] ? GRReg_18 : _GEN_17; // @[GRReg.scala 24:{24,24}]
  wire [63:0] _GEN_19 = 6'h13 == io_rj_addr[5:0] ? GRReg_19 : _GEN_18; // @[GRReg.scala 24:{24,24}]
  wire [63:0] _GEN_20 = 6'h14 == io_rj_addr[5:0] ? GRReg_20 : _GEN_19; // @[GRReg.scala 24:{24,24}]
  wire [63:0] _GEN_21 = 6'h15 == io_rj_addr[5:0] ? GRReg_21 : _GEN_20; // @[GRReg.scala 24:{24,24}]
  wire [63:0] _GEN_22 = 6'h16 == io_rj_addr[5:0] ? GRReg_22 : _GEN_21; // @[GRReg.scala 24:{24,24}]
  wire [63:0] _GEN_23 = 6'h17 == io_rj_addr[5:0] ? GRReg_23 : _GEN_22; // @[GRReg.scala 24:{24,24}]
  wire [63:0] _GEN_24 = 6'h18 == io_rj_addr[5:0] ? GRReg_24 : _GEN_23; // @[GRReg.scala 24:{24,24}]
  wire [63:0] _GEN_25 = 6'h19 == io_rj_addr[5:0] ? GRReg_25 : _GEN_24; // @[GRReg.scala 24:{24,24}]
  wire [63:0] _GEN_26 = 6'h1a == io_rj_addr[5:0] ? GRReg_26 : _GEN_25; // @[GRReg.scala 24:{24,24}]
  wire [63:0] _GEN_27 = 6'h1b == io_rj_addr[5:0] ? GRReg_27 : _GEN_26; // @[GRReg.scala 24:{24,24}]
  wire [63:0] _GEN_28 = 6'h1c == io_rj_addr[5:0] ? GRReg_28 : _GEN_27; // @[GRReg.scala 24:{24,24}]
  wire [63:0] _GEN_29 = 6'h1d == io_rj_addr[5:0] ? GRReg_29 : _GEN_28; // @[GRReg.scala 24:{24,24}]
  wire [63:0] _GEN_30 = 6'h1e == io_rj_addr[5:0] ? GRReg_30 : _GEN_29; // @[GRReg.scala 24:{24,24}]
  wire [63:0] _GEN_31 = 6'h1f == io_rj_addr[5:0] ? GRReg_31 : _GEN_30; // @[GRReg.scala 24:{24,24}]
  wire [63:0] _GEN_32 = 6'h20 == io_rj_addr[5:0] ? GRReg_32 : _GEN_31; // @[GRReg.scala 24:{24,24}]
  wire [63:0] _GEN_33 = 6'h21 == io_rj_addr[5:0] ? GRReg_33 : _GEN_32; // @[GRReg.scala 24:{24,24}]
  wire [63:0] _GEN_34 = 6'h22 == io_rj_addr[5:0] ? GRReg_34 : _GEN_33; // @[GRReg.scala 24:{24,24}]
  wire [63:0] _GEN_35 = 6'h23 == io_rj_addr[5:0] ? GRReg_35 : _GEN_34; // @[GRReg.scala 24:{24,24}]
  wire [63:0] _GEN_36 = 6'h24 == io_rj_addr[5:0] ? GRReg_36 : _GEN_35; // @[GRReg.scala 24:{24,24}]
  wire [63:0] _GEN_37 = 6'h25 == io_rj_addr[5:0] ? GRReg_37 : _GEN_36; // @[GRReg.scala 24:{24,24}]
  wire [63:0] _GEN_38 = 6'h26 == io_rj_addr[5:0] ? GRReg_38 : _GEN_37; // @[GRReg.scala 24:{24,24}]
  wire [63:0] _GEN_39 = 6'h27 == io_rj_addr[5:0] ? GRReg_39 : _GEN_38; // @[GRReg.scala 24:{24,24}]
  wire [63:0] _GEN_40 = 6'h28 == io_rj_addr[5:0] ? GRReg_40 : _GEN_39; // @[GRReg.scala 24:{24,24}]
  wire [63:0] _GEN_41 = 6'h29 == io_rj_addr[5:0] ? GRReg_41 : _GEN_40; // @[GRReg.scala 24:{24,24}]
  wire [63:0] _GEN_42 = 6'h2a == io_rj_addr[5:0] ? GRReg_42 : _GEN_41; // @[GRReg.scala 24:{24,24}]
  wire [63:0] _GEN_43 = 6'h2b == io_rj_addr[5:0] ? GRReg_43 : _GEN_42; // @[GRReg.scala 24:{24,24}]
  wire [63:0] _GEN_44 = 6'h2c == io_rj_addr[5:0] ? GRReg_44 : _GEN_43; // @[GRReg.scala 24:{24,24}]
  wire [63:0] _GEN_45 = 6'h2d == io_rj_addr[5:0] ? GRReg_45 : _GEN_44; // @[GRReg.scala 24:{24,24}]
  wire [63:0] _GEN_46 = 6'h2e == io_rj_addr[5:0] ? GRReg_46 : _GEN_45; // @[GRReg.scala 24:{24,24}]
  wire [63:0] _GEN_47 = 6'h2f == io_rj_addr[5:0] ? GRReg_47 : _GEN_46; // @[GRReg.scala 24:{24,24}]
  wire [63:0] _GEN_48 = 6'h30 == io_rj_addr[5:0] ? GRReg_48 : _GEN_47; // @[GRReg.scala 24:{24,24}]
  wire [63:0] _GEN_49 = 6'h31 == io_rj_addr[5:0] ? GRReg_49 : _GEN_48; // @[GRReg.scala 24:{24,24}]
  wire [63:0] _GEN_50 = 6'h32 == io_rj_addr[5:0] ? GRReg_50 : _GEN_49; // @[GRReg.scala 24:{24,24}]
  wire [63:0] _GEN_51 = 6'h33 == io_rj_addr[5:0] ? GRReg_51 : _GEN_50; // @[GRReg.scala 24:{24,24}]
  wire [63:0] _GEN_52 = 6'h34 == io_rj_addr[5:0] ? GRReg_52 : _GEN_51; // @[GRReg.scala 24:{24,24}]
  wire [63:0] _GEN_53 = 6'h35 == io_rj_addr[5:0] ? GRReg_53 : _GEN_52; // @[GRReg.scala 24:{24,24}]
  wire [63:0] _GEN_54 = 6'h36 == io_rj_addr[5:0] ? GRReg_54 : _GEN_53; // @[GRReg.scala 24:{24,24}]
  wire [63:0] _GEN_55 = 6'h37 == io_rj_addr[5:0] ? GRReg_55 : _GEN_54; // @[GRReg.scala 24:{24,24}]
  wire [63:0] _GEN_56 = 6'h38 == io_rj_addr[5:0] ? GRReg_56 : _GEN_55; // @[GRReg.scala 24:{24,24}]
  wire [63:0] _GEN_57 = 6'h39 == io_rj_addr[5:0] ? GRReg_57 : _GEN_56; // @[GRReg.scala 24:{24,24}]
  wire [63:0] _GEN_58 = 6'h3a == io_rj_addr[5:0] ? GRReg_58 : _GEN_57; // @[GRReg.scala 24:{24,24}]
  wire [63:0] _GEN_59 = 6'h3b == io_rj_addr[5:0] ? GRReg_59 : _GEN_58; // @[GRReg.scala 24:{24,24}]
  wire [63:0] _GEN_60 = 6'h3c == io_rj_addr[5:0] ? GRReg_60 : _GEN_59; // @[GRReg.scala 24:{24,24}]
  wire [63:0] _GEN_61 = 6'h3d == io_rj_addr[5:0] ? GRReg_61 : _GEN_60; // @[GRReg.scala 24:{24,24}]
  wire [63:0] _GEN_62 = 6'h3e == io_rj_addr[5:0] ? GRReg_62 : _GEN_61; // @[GRReg.scala 24:{24,24}]
  wire [63:0] _GEN_65 = 6'h1 == io_rk_addr[5:0] ? GRReg_1 : GRReg_0; // @[GRReg.scala 25:{24,24}]
  wire [63:0] _GEN_66 = 6'h2 == io_rk_addr[5:0] ? GRReg_2 : _GEN_65; // @[GRReg.scala 25:{24,24}]
  wire [63:0] _GEN_67 = 6'h3 == io_rk_addr[5:0] ? GRReg_3 : _GEN_66; // @[GRReg.scala 25:{24,24}]
  wire [63:0] _GEN_68 = 6'h4 == io_rk_addr[5:0] ? GRReg_4 : _GEN_67; // @[GRReg.scala 25:{24,24}]
  wire [63:0] _GEN_69 = 6'h5 == io_rk_addr[5:0] ? GRReg_5 : _GEN_68; // @[GRReg.scala 25:{24,24}]
  wire [63:0] _GEN_70 = 6'h6 == io_rk_addr[5:0] ? GRReg_6 : _GEN_69; // @[GRReg.scala 25:{24,24}]
  wire [63:0] _GEN_71 = 6'h7 == io_rk_addr[5:0] ? GRReg_7 : _GEN_70; // @[GRReg.scala 25:{24,24}]
  wire [63:0] _GEN_72 = 6'h8 == io_rk_addr[5:0] ? GRReg_8 : _GEN_71; // @[GRReg.scala 25:{24,24}]
  wire [63:0] _GEN_73 = 6'h9 == io_rk_addr[5:0] ? GRReg_9 : _GEN_72; // @[GRReg.scala 25:{24,24}]
  wire [63:0] _GEN_74 = 6'ha == io_rk_addr[5:0] ? GRReg_10 : _GEN_73; // @[GRReg.scala 25:{24,24}]
  wire [63:0] _GEN_75 = 6'hb == io_rk_addr[5:0] ? GRReg_11 : _GEN_74; // @[GRReg.scala 25:{24,24}]
  wire [63:0] _GEN_76 = 6'hc == io_rk_addr[5:0] ? GRReg_12 : _GEN_75; // @[GRReg.scala 25:{24,24}]
  wire [63:0] _GEN_77 = 6'hd == io_rk_addr[5:0] ? GRReg_13 : _GEN_76; // @[GRReg.scala 25:{24,24}]
  wire [63:0] _GEN_78 = 6'he == io_rk_addr[5:0] ? GRReg_14 : _GEN_77; // @[GRReg.scala 25:{24,24}]
  wire [63:0] _GEN_79 = 6'hf == io_rk_addr[5:0] ? GRReg_15 : _GEN_78; // @[GRReg.scala 25:{24,24}]
  wire [63:0] _GEN_80 = 6'h10 == io_rk_addr[5:0] ? GRReg_16 : _GEN_79; // @[GRReg.scala 25:{24,24}]
  wire [63:0] _GEN_81 = 6'h11 == io_rk_addr[5:0] ? GRReg_17 : _GEN_80; // @[GRReg.scala 25:{24,24}]
  wire [63:0] _GEN_82 = 6'h12 == io_rk_addr[5:0] ? GRReg_18 : _GEN_81; // @[GRReg.scala 25:{24,24}]
  wire [63:0] _GEN_83 = 6'h13 == io_rk_addr[5:0] ? GRReg_19 : _GEN_82; // @[GRReg.scala 25:{24,24}]
  wire [63:0] _GEN_84 = 6'h14 == io_rk_addr[5:0] ? GRReg_20 : _GEN_83; // @[GRReg.scala 25:{24,24}]
  wire [63:0] _GEN_85 = 6'h15 == io_rk_addr[5:0] ? GRReg_21 : _GEN_84; // @[GRReg.scala 25:{24,24}]
  wire [63:0] _GEN_86 = 6'h16 == io_rk_addr[5:0] ? GRReg_22 : _GEN_85; // @[GRReg.scala 25:{24,24}]
  wire [63:0] _GEN_87 = 6'h17 == io_rk_addr[5:0] ? GRReg_23 : _GEN_86; // @[GRReg.scala 25:{24,24}]
  wire [63:0] _GEN_88 = 6'h18 == io_rk_addr[5:0] ? GRReg_24 : _GEN_87; // @[GRReg.scala 25:{24,24}]
  wire [63:0] _GEN_89 = 6'h19 == io_rk_addr[5:0] ? GRReg_25 : _GEN_88; // @[GRReg.scala 25:{24,24}]
  wire [63:0] _GEN_90 = 6'h1a == io_rk_addr[5:0] ? GRReg_26 : _GEN_89; // @[GRReg.scala 25:{24,24}]
  wire [63:0] _GEN_91 = 6'h1b == io_rk_addr[5:0] ? GRReg_27 : _GEN_90; // @[GRReg.scala 25:{24,24}]
  wire [63:0] _GEN_92 = 6'h1c == io_rk_addr[5:0] ? GRReg_28 : _GEN_91; // @[GRReg.scala 25:{24,24}]
  wire [63:0] _GEN_93 = 6'h1d == io_rk_addr[5:0] ? GRReg_29 : _GEN_92; // @[GRReg.scala 25:{24,24}]
  wire [63:0] _GEN_94 = 6'h1e == io_rk_addr[5:0] ? GRReg_30 : _GEN_93; // @[GRReg.scala 25:{24,24}]
  wire [63:0] _GEN_95 = 6'h1f == io_rk_addr[5:0] ? GRReg_31 : _GEN_94; // @[GRReg.scala 25:{24,24}]
  wire [63:0] _GEN_96 = 6'h20 == io_rk_addr[5:0] ? GRReg_32 : _GEN_95; // @[GRReg.scala 25:{24,24}]
  wire [63:0] _GEN_97 = 6'h21 == io_rk_addr[5:0] ? GRReg_33 : _GEN_96; // @[GRReg.scala 25:{24,24}]
  wire [63:0] _GEN_98 = 6'h22 == io_rk_addr[5:0] ? GRReg_34 : _GEN_97; // @[GRReg.scala 25:{24,24}]
  wire [63:0] _GEN_99 = 6'h23 == io_rk_addr[5:0] ? GRReg_35 : _GEN_98; // @[GRReg.scala 25:{24,24}]
  wire [63:0] _GEN_100 = 6'h24 == io_rk_addr[5:0] ? GRReg_36 : _GEN_99; // @[GRReg.scala 25:{24,24}]
  wire [63:0] _GEN_101 = 6'h25 == io_rk_addr[5:0] ? GRReg_37 : _GEN_100; // @[GRReg.scala 25:{24,24}]
  wire [63:0] _GEN_102 = 6'h26 == io_rk_addr[5:0] ? GRReg_38 : _GEN_101; // @[GRReg.scala 25:{24,24}]
  wire [63:0] _GEN_103 = 6'h27 == io_rk_addr[5:0] ? GRReg_39 : _GEN_102; // @[GRReg.scala 25:{24,24}]
  wire [63:0] _GEN_104 = 6'h28 == io_rk_addr[5:0] ? GRReg_40 : _GEN_103; // @[GRReg.scala 25:{24,24}]
  wire [63:0] _GEN_105 = 6'h29 == io_rk_addr[5:0] ? GRReg_41 : _GEN_104; // @[GRReg.scala 25:{24,24}]
  wire [63:0] _GEN_106 = 6'h2a == io_rk_addr[5:0] ? GRReg_42 : _GEN_105; // @[GRReg.scala 25:{24,24}]
  wire [63:0] _GEN_107 = 6'h2b == io_rk_addr[5:0] ? GRReg_43 : _GEN_106; // @[GRReg.scala 25:{24,24}]
  wire [63:0] _GEN_108 = 6'h2c == io_rk_addr[5:0] ? GRReg_44 : _GEN_107; // @[GRReg.scala 25:{24,24}]
  wire [63:0] _GEN_109 = 6'h2d == io_rk_addr[5:0] ? GRReg_45 : _GEN_108; // @[GRReg.scala 25:{24,24}]
  wire [63:0] _GEN_110 = 6'h2e == io_rk_addr[5:0] ? GRReg_46 : _GEN_109; // @[GRReg.scala 25:{24,24}]
  wire [63:0] _GEN_111 = 6'h2f == io_rk_addr[5:0] ? GRReg_47 : _GEN_110; // @[GRReg.scala 25:{24,24}]
  wire [63:0] _GEN_112 = 6'h30 == io_rk_addr[5:0] ? GRReg_48 : _GEN_111; // @[GRReg.scala 25:{24,24}]
  wire [63:0] _GEN_113 = 6'h31 == io_rk_addr[5:0] ? GRReg_49 : _GEN_112; // @[GRReg.scala 25:{24,24}]
  wire [63:0] _GEN_114 = 6'h32 == io_rk_addr[5:0] ? GRReg_50 : _GEN_113; // @[GRReg.scala 25:{24,24}]
  wire [63:0] _GEN_115 = 6'h33 == io_rk_addr[5:0] ? GRReg_51 : _GEN_114; // @[GRReg.scala 25:{24,24}]
  wire [63:0] _GEN_116 = 6'h34 == io_rk_addr[5:0] ? GRReg_52 : _GEN_115; // @[GRReg.scala 25:{24,24}]
  wire [63:0] _GEN_117 = 6'h35 == io_rk_addr[5:0] ? GRReg_53 : _GEN_116; // @[GRReg.scala 25:{24,24}]
  wire [63:0] _GEN_118 = 6'h36 == io_rk_addr[5:0] ? GRReg_54 : _GEN_117; // @[GRReg.scala 25:{24,24}]
  wire [63:0] _GEN_119 = 6'h37 == io_rk_addr[5:0] ? GRReg_55 : _GEN_118; // @[GRReg.scala 25:{24,24}]
  wire [63:0] _GEN_120 = 6'h38 == io_rk_addr[5:0] ? GRReg_56 : _GEN_119; // @[GRReg.scala 25:{24,24}]
  wire [63:0] _GEN_121 = 6'h39 == io_rk_addr[5:0] ? GRReg_57 : _GEN_120; // @[GRReg.scala 25:{24,24}]
  wire [63:0] _GEN_122 = 6'h3a == io_rk_addr[5:0] ? GRReg_58 : _GEN_121; // @[GRReg.scala 25:{24,24}]
  wire [63:0] _GEN_123 = 6'h3b == io_rk_addr[5:0] ? GRReg_59 : _GEN_122; // @[GRReg.scala 25:{24,24}]
  wire [63:0] _GEN_124 = 6'h3c == io_rk_addr[5:0] ? GRReg_60 : _GEN_123; // @[GRReg.scala 25:{24,24}]
  wire [63:0] _GEN_125 = 6'h3d == io_rk_addr[5:0] ? GRReg_61 : _GEN_124; // @[GRReg.scala 25:{24,24}]
  wire [63:0] _GEN_126 = 6'h3e == io_rk_addr[5:0] ? GRReg_62 : _GEN_125; // @[GRReg.scala 25:{24,24}]
  wire [63:0] _GEN_129 = 6'h1 == io_rd_addr[5:0] ? GRReg_1 : GRReg_0; // @[GRReg.scala 26:{27,27}]
  wire [63:0] _GEN_130 = 6'h2 == io_rd_addr[5:0] ? GRReg_2 : _GEN_129; // @[GRReg.scala 26:{27,27}]
  wire [63:0] _GEN_131 = 6'h3 == io_rd_addr[5:0] ? GRReg_3 : _GEN_130; // @[GRReg.scala 26:{27,27}]
  wire [63:0] _GEN_132 = 6'h4 == io_rd_addr[5:0] ? GRReg_4 : _GEN_131; // @[GRReg.scala 26:{27,27}]
  wire [63:0] _GEN_133 = 6'h5 == io_rd_addr[5:0] ? GRReg_5 : _GEN_132; // @[GRReg.scala 26:{27,27}]
  wire [63:0] _GEN_134 = 6'h6 == io_rd_addr[5:0] ? GRReg_6 : _GEN_133; // @[GRReg.scala 26:{27,27}]
  wire [63:0] _GEN_135 = 6'h7 == io_rd_addr[5:0] ? GRReg_7 : _GEN_134; // @[GRReg.scala 26:{27,27}]
  wire [63:0] _GEN_136 = 6'h8 == io_rd_addr[5:0] ? GRReg_8 : _GEN_135; // @[GRReg.scala 26:{27,27}]
  wire [63:0] _GEN_137 = 6'h9 == io_rd_addr[5:0] ? GRReg_9 : _GEN_136; // @[GRReg.scala 26:{27,27}]
  wire [63:0] _GEN_138 = 6'ha == io_rd_addr[5:0] ? GRReg_10 : _GEN_137; // @[GRReg.scala 26:{27,27}]
  wire [63:0] _GEN_139 = 6'hb == io_rd_addr[5:0] ? GRReg_11 : _GEN_138; // @[GRReg.scala 26:{27,27}]
  wire [63:0] _GEN_140 = 6'hc == io_rd_addr[5:0] ? GRReg_12 : _GEN_139; // @[GRReg.scala 26:{27,27}]
  wire [63:0] _GEN_141 = 6'hd == io_rd_addr[5:0] ? GRReg_13 : _GEN_140; // @[GRReg.scala 26:{27,27}]
  wire [63:0] _GEN_142 = 6'he == io_rd_addr[5:0] ? GRReg_14 : _GEN_141; // @[GRReg.scala 26:{27,27}]
  wire [63:0] _GEN_143 = 6'hf == io_rd_addr[5:0] ? GRReg_15 : _GEN_142; // @[GRReg.scala 26:{27,27}]
  wire [63:0] _GEN_144 = 6'h10 == io_rd_addr[5:0] ? GRReg_16 : _GEN_143; // @[GRReg.scala 26:{27,27}]
  wire [63:0] _GEN_145 = 6'h11 == io_rd_addr[5:0] ? GRReg_17 : _GEN_144; // @[GRReg.scala 26:{27,27}]
  wire [63:0] _GEN_146 = 6'h12 == io_rd_addr[5:0] ? GRReg_18 : _GEN_145; // @[GRReg.scala 26:{27,27}]
  wire [63:0] _GEN_147 = 6'h13 == io_rd_addr[5:0] ? GRReg_19 : _GEN_146; // @[GRReg.scala 26:{27,27}]
  wire [63:0] _GEN_148 = 6'h14 == io_rd_addr[5:0] ? GRReg_20 : _GEN_147; // @[GRReg.scala 26:{27,27}]
  wire [63:0] _GEN_149 = 6'h15 == io_rd_addr[5:0] ? GRReg_21 : _GEN_148; // @[GRReg.scala 26:{27,27}]
  wire [63:0] _GEN_150 = 6'h16 == io_rd_addr[5:0] ? GRReg_22 : _GEN_149; // @[GRReg.scala 26:{27,27}]
  wire [63:0] _GEN_151 = 6'h17 == io_rd_addr[5:0] ? GRReg_23 : _GEN_150; // @[GRReg.scala 26:{27,27}]
  wire [63:0] _GEN_152 = 6'h18 == io_rd_addr[5:0] ? GRReg_24 : _GEN_151; // @[GRReg.scala 26:{27,27}]
  wire [63:0] _GEN_153 = 6'h19 == io_rd_addr[5:0] ? GRReg_25 : _GEN_152; // @[GRReg.scala 26:{27,27}]
  wire [63:0] _GEN_154 = 6'h1a == io_rd_addr[5:0] ? GRReg_26 : _GEN_153; // @[GRReg.scala 26:{27,27}]
  wire [63:0] _GEN_155 = 6'h1b == io_rd_addr[5:0] ? GRReg_27 : _GEN_154; // @[GRReg.scala 26:{27,27}]
  wire [63:0] _GEN_156 = 6'h1c == io_rd_addr[5:0] ? GRReg_28 : _GEN_155; // @[GRReg.scala 26:{27,27}]
  wire [63:0] _GEN_157 = 6'h1d == io_rd_addr[5:0] ? GRReg_29 : _GEN_156; // @[GRReg.scala 26:{27,27}]
  wire [63:0] _GEN_158 = 6'h1e == io_rd_addr[5:0] ? GRReg_30 : _GEN_157; // @[GRReg.scala 26:{27,27}]
  wire [63:0] _GEN_159 = 6'h1f == io_rd_addr[5:0] ? GRReg_31 : _GEN_158; // @[GRReg.scala 26:{27,27}]
  wire [63:0] _GEN_160 = 6'h20 == io_rd_addr[5:0] ? GRReg_32 : _GEN_159; // @[GRReg.scala 26:{27,27}]
  wire [63:0] _GEN_161 = 6'h21 == io_rd_addr[5:0] ? GRReg_33 : _GEN_160; // @[GRReg.scala 26:{27,27}]
  wire [63:0] _GEN_162 = 6'h22 == io_rd_addr[5:0] ? GRReg_34 : _GEN_161; // @[GRReg.scala 26:{27,27}]
  wire [63:0] _GEN_163 = 6'h23 == io_rd_addr[5:0] ? GRReg_35 : _GEN_162; // @[GRReg.scala 26:{27,27}]
  wire [63:0] _GEN_164 = 6'h24 == io_rd_addr[5:0] ? GRReg_36 : _GEN_163; // @[GRReg.scala 26:{27,27}]
  wire [63:0] _GEN_165 = 6'h25 == io_rd_addr[5:0] ? GRReg_37 : _GEN_164; // @[GRReg.scala 26:{27,27}]
  wire [63:0] _GEN_166 = 6'h26 == io_rd_addr[5:0] ? GRReg_38 : _GEN_165; // @[GRReg.scala 26:{27,27}]
  wire [63:0] _GEN_167 = 6'h27 == io_rd_addr[5:0] ? GRReg_39 : _GEN_166; // @[GRReg.scala 26:{27,27}]
  wire [63:0] _GEN_168 = 6'h28 == io_rd_addr[5:0] ? GRReg_40 : _GEN_167; // @[GRReg.scala 26:{27,27}]
  wire [63:0] _GEN_169 = 6'h29 == io_rd_addr[5:0] ? GRReg_41 : _GEN_168; // @[GRReg.scala 26:{27,27}]
  wire [63:0] _GEN_170 = 6'h2a == io_rd_addr[5:0] ? GRReg_42 : _GEN_169; // @[GRReg.scala 26:{27,27}]
  wire [63:0] _GEN_171 = 6'h2b == io_rd_addr[5:0] ? GRReg_43 : _GEN_170; // @[GRReg.scala 26:{27,27}]
  wire [63:0] _GEN_172 = 6'h2c == io_rd_addr[5:0] ? GRReg_44 : _GEN_171; // @[GRReg.scala 26:{27,27}]
  wire [63:0] _GEN_173 = 6'h2d == io_rd_addr[5:0] ? GRReg_45 : _GEN_172; // @[GRReg.scala 26:{27,27}]
  wire [63:0] _GEN_174 = 6'h2e == io_rd_addr[5:0] ? GRReg_46 : _GEN_173; // @[GRReg.scala 26:{27,27}]
  wire [63:0] _GEN_175 = 6'h2f == io_rd_addr[5:0] ? GRReg_47 : _GEN_174; // @[GRReg.scala 26:{27,27}]
  wire [63:0] _GEN_176 = 6'h30 == io_rd_addr[5:0] ? GRReg_48 : _GEN_175; // @[GRReg.scala 26:{27,27}]
  wire [63:0] _GEN_177 = 6'h31 == io_rd_addr[5:0] ? GRReg_49 : _GEN_176; // @[GRReg.scala 26:{27,27}]
  wire [63:0] _GEN_178 = 6'h32 == io_rd_addr[5:0] ? GRReg_50 : _GEN_177; // @[GRReg.scala 26:{27,27}]
  wire [63:0] _GEN_179 = 6'h33 == io_rd_addr[5:0] ? GRReg_51 : _GEN_178; // @[GRReg.scala 26:{27,27}]
  wire [63:0] _GEN_180 = 6'h34 == io_rd_addr[5:0] ? GRReg_52 : _GEN_179; // @[GRReg.scala 26:{27,27}]
  wire [63:0] _GEN_181 = 6'h35 == io_rd_addr[5:0] ? GRReg_53 : _GEN_180; // @[GRReg.scala 26:{27,27}]
  wire [63:0] _GEN_182 = 6'h36 == io_rd_addr[5:0] ? GRReg_54 : _GEN_181; // @[GRReg.scala 26:{27,27}]
  wire [63:0] _GEN_183 = 6'h37 == io_rd_addr[5:0] ? GRReg_55 : _GEN_182; // @[GRReg.scala 26:{27,27}]
  wire [63:0] _GEN_184 = 6'h38 == io_rd_addr[5:0] ? GRReg_56 : _GEN_183; // @[GRReg.scala 26:{27,27}]
  wire [63:0] _GEN_185 = 6'h39 == io_rd_addr[5:0] ? GRReg_57 : _GEN_184; // @[GRReg.scala 26:{27,27}]
  wire [63:0] _GEN_186 = 6'h3a == io_rd_addr[5:0] ? GRReg_58 : _GEN_185; // @[GRReg.scala 26:{27,27}]
  wire [63:0] _GEN_187 = 6'h3b == io_rd_addr[5:0] ? GRReg_59 : _GEN_186; // @[GRReg.scala 26:{27,27}]
  wire [63:0] _GEN_188 = 6'h3c == io_rd_addr[5:0] ? GRReg_60 : _GEN_187; // @[GRReg.scala 26:{27,27}]
  wire [63:0] _GEN_189 = 6'h3d == io_rd_addr[5:0] ? GRReg_61 : _GEN_188; // @[GRReg.scala 26:{27,27}]
  wire [63:0] _GEN_190 = 6'h3e == io_rd_addr[5:0] ? GRReg_62 : _GEN_189; // @[GRReg.scala 26:{27,27}]
  assign io_ALU_GRReg_IO_rj = 6'h3f == io_rj_addr[5:0] ? GRReg_63 : _GEN_62; // @[GRReg.scala 24:{24,24}]
  assign io_ALU_GRReg_IO_rk = 6'h3f == io_rk_addr[5:0] ? GRReg_63 : _GEN_126; // @[GRReg.scala 25:{24,24}]
  assign io_ALU_GRReg_IO_rd_in = 6'h3f == io_rd_addr[5:0] ? GRReg_63 : _GEN_190; // @[GRReg.scala 26:{27,27}]
  always @(posedge clock) begin
    if (reset) begin // @[GRReg.scala 22:24]
      GRReg_0 <= 64'h0; // @[GRReg.scala 22:24]
    end else if (6'h0 == io_rd_addr[5:0]) begin // @[GRReg.scala 28:23]
      GRReg_0 <= io_ALU_GRReg_IO_rd; // @[GRReg.scala 28:23]
    end
    if (reset) begin // @[GRReg.scala 22:24]
      GRReg_1 <= 64'h0; // @[GRReg.scala 22:24]
    end else if (6'h1 == io_rd_addr[5:0]) begin // @[GRReg.scala 28:23]
      GRReg_1 <= io_ALU_GRReg_IO_rd; // @[GRReg.scala 28:23]
    end
    if (reset) begin // @[GRReg.scala 22:24]
      GRReg_2 <= 64'h0; // @[GRReg.scala 22:24]
    end else if (6'h2 == io_rd_addr[5:0]) begin // @[GRReg.scala 28:23]
      GRReg_2 <= io_ALU_GRReg_IO_rd; // @[GRReg.scala 28:23]
    end
    if (reset) begin // @[GRReg.scala 22:24]
      GRReg_3 <= 64'h0; // @[GRReg.scala 22:24]
    end else if (6'h3 == io_rd_addr[5:0]) begin // @[GRReg.scala 28:23]
      GRReg_3 <= io_ALU_GRReg_IO_rd; // @[GRReg.scala 28:23]
    end
    if (reset) begin // @[GRReg.scala 22:24]
      GRReg_4 <= 64'h0; // @[GRReg.scala 22:24]
    end else if (6'h4 == io_rd_addr[5:0]) begin // @[GRReg.scala 28:23]
      GRReg_4 <= io_ALU_GRReg_IO_rd; // @[GRReg.scala 28:23]
    end
    if (reset) begin // @[GRReg.scala 22:24]
      GRReg_5 <= 64'h0; // @[GRReg.scala 22:24]
    end else if (6'h5 == io_rd_addr[5:0]) begin // @[GRReg.scala 28:23]
      GRReg_5 <= io_ALU_GRReg_IO_rd; // @[GRReg.scala 28:23]
    end
    if (reset) begin // @[GRReg.scala 22:24]
      GRReg_6 <= 64'h0; // @[GRReg.scala 22:24]
    end else if (6'h6 == io_rd_addr[5:0]) begin // @[GRReg.scala 28:23]
      GRReg_6 <= io_ALU_GRReg_IO_rd; // @[GRReg.scala 28:23]
    end
    if (reset) begin // @[GRReg.scala 22:24]
      GRReg_7 <= 64'h0; // @[GRReg.scala 22:24]
    end else if (6'h7 == io_rd_addr[5:0]) begin // @[GRReg.scala 28:23]
      GRReg_7 <= io_ALU_GRReg_IO_rd; // @[GRReg.scala 28:23]
    end
    if (reset) begin // @[GRReg.scala 22:24]
      GRReg_8 <= 64'h0; // @[GRReg.scala 22:24]
    end else if (6'h8 == io_rd_addr[5:0]) begin // @[GRReg.scala 28:23]
      GRReg_8 <= io_ALU_GRReg_IO_rd; // @[GRReg.scala 28:23]
    end
    if (reset) begin // @[GRReg.scala 22:24]
      GRReg_9 <= 64'h0; // @[GRReg.scala 22:24]
    end else if (6'h9 == io_rd_addr[5:0]) begin // @[GRReg.scala 28:23]
      GRReg_9 <= io_ALU_GRReg_IO_rd; // @[GRReg.scala 28:23]
    end
    if (reset) begin // @[GRReg.scala 22:24]
      GRReg_10 <= 64'h0; // @[GRReg.scala 22:24]
    end else if (6'ha == io_rd_addr[5:0]) begin // @[GRReg.scala 28:23]
      GRReg_10 <= io_ALU_GRReg_IO_rd; // @[GRReg.scala 28:23]
    end
    if (reset) begin // @[GRReg.scala 22:24]
      GRReg_11 <= 64'h0; // @[GRReg.scala 22:24]
    end else if (6'hb == io_rd_addr[5:0]) begin // @[GRReg.scala 28:23]
      GRReg_11 <= io_ALU_GRReg_IO_rd; // @[GRReg.scala 28:23]
    end
    if (reset) begin // @[GRReg.scala 22:24]
      GRReg_12 <= 64'h0; // @[GRReg.scala 22:24]
    end else if (6'hc == io_rd_addr[5:0]) begin // @[GRReg.scala 28:23]
      GRReg_12 <= io_ALU_GRReg_IO_rd; // @[GRReg.scala 28:23]
    end
    if (reset) begin // @[GRReg.scala 22:24]
      GRReg_13 <= 64'h0; // @[GRReg.scala 22:24]
    end else if (6'hd == io_rd_addr[5:0]) begin // @[GRReg.scala 28:23]
      GRReg_13 <= io_ALU_GRReg_IO_rd; // @[GRReg.scala 28:23]
    end
    if (reset) begin // @[GRReg.scala 22:24]
      GRReg_14 <= 64'h0; // @[GRReg.scala 22:24]
    end else if (6'he == io_rd_addr[5:0]) begin // @[GRReg.scala 28:23]
      GRReg_14 <= io_ALU_GRReg_IO_rd; // @[GRReg.scala 28:23]
    end
    if (reset) begin // @[GRReg.scala 22:24]
      GRReg_15 <= 64'h0; // @[GRReg.scala 22:24]
    end else if (6'hf == io_rd_addr[5:0]) begin // @[GRReg.scala 28:23]
      GRReg_15 <= io_ALU_GRReg_IO_rd; // @[GRReg.scala 28:23]
    end
    if (reset) begin // @[GRReg.scala 22:24]
      GRReg_16 <= 64'h0; // @[GRReg.scala 22:24]
    end else if (6'h10 == io_rd_addr[5:0]) begin // @[GRReg.scala 28:23]
      GRReg_16 <= io_ALU_GRReg_IO_rd; // @[GRReg.scala 28:23]
    end
    if (reset) begin // @[GRReg.scala 22:24]
      GRReg_17 <= 64'h0; // @[GRReg.scala 22:24]
    end else if (6'h11 == io_rd_addr[5:0]) begin // @[GRReg.scala 28:23]
      GRReg_17 <= io_ALU_GRReg_IO_rd; // @[GRReg.scala 28:23]
    end
    if (reset) begin // @[GRReg.scala 22:24]
      GRReg_18 <= 64'h0; // @[GRReg.scala 22:24]
    end else if (6'h12 == io_rd_addr[5:0]) begin // @[GRReg.scala 28:23]
      GRReg_18 <= io_ALU_GRReg_IO_rd; // @[GRReg.scala 28:23]
    end
    if (reset) begin // @[GRReg.scala 22:24]
      GRReg_19 <= 64'h0; // @[GRReg.scala 22:24]
    end else if (6'h13 == io_rd_addr[5:0]) begin // @[GRReg.scala 28:23]
      GRReg_19 <= io_ALU_GRReg_IO_rd; // @[GRReg.scala 28:23]
    end
    if (reset) begin // @[GRReg.scala 22:24]
      GRReg_20 <= 64'h0; // @[GRReg.scala 22:24]
    end else if (6'h14 == io_rd_addr[5:0]) begin // @[GRReg.scala 28:23]
      GRReg_20 <= io_ALU_GRReg_IO_rd; // @[GRReg.scala 28:23]
    end
    if (reset) begin // @[GRReg.scala 22:24]
      GRReg_21 <= 64'h0; // @[GRReg.scala 22:24]
    end else if (6'h15 == io_rd_addr[5:0]) begin // @[GRReg.scala 28:23]
      GRReg_21 <= io_ALU_GRReg_IO_rd; // @[GRReg.scala 28:23]
    end
    if (reset) begin // @[GRReg.scala 22:24]
      GRReg_22 <= 64'h0; // @[GRReg.scala 22:24]
    end else if (6'h16 == io_rd_addr[5:0]) begin // @[GRReg.scala 28:23]
      GRReg_22 <= io_ALU_GRReg_IO_rd; // @[GRReg.scala 28:23]
    end
    if (reset) begin // @[GRReg.scala 22:24]
      GRReg_23 <= 64'h0; // @[GRReg.scala 22:24]
    end else if (6'h17 == io_rd_addr[5:0]) begin // @[GRReg.scala 28:23]
      GRReg_23 <= io_ALU_GRReg_IO_rd; // @[GRReg.scala 28:23]
    end
    if (reset) begin // @[GRReg.scala 22:24]
      GRReg_24 <= 64'h0; // @[GRReg.scala 22:24]
    end else if (6'h18 == io_rd_addr[5:0]) begin // @[GRReg.scala 28:23]
      GRReg_24 <= io_ALU_GRReg_IO_rd; // @[GRReg.scala 28:23]
    end
    if (reset) begin // @[GRReg.scala 22:24]
      GRReg_25 <= 64'h0; // @[GRReg.scala 22:24]
    end else if (6'h19 == io_rd_addr[5:0]) begin // @[GRReg.scala 28:23]
      GRReg_25 <= io_ALU_GRReg_IO_rd; // @[GRReg.scala 28:23]
    end
    if (reset) begin // @[GRReg.scala 22:24]
      GRReg_26 <= 64'h0; // @[GRReg.scala 22:24]
    end else if (6'h1a == io_rd_addr[5:0]) begin // @[GRReg.scala 28:23]
      GRReg_26 <= io_ALU_GRReg_IO_rd; // @[GRReg.scala 28:23]
    end
    if (reset) begin // @[GRReg.scala 22:24]
      GRReg_27 <= 64'h0; // @[GRReg.scala 22:24]
    end else if (6'h1b == io_rd_addr[5:0]) begin // @[GRReg.scala 28:23]
      GRReg_27 <= io_ALU_GRReg_IO_rd; // @[GRReg.scala 28:23]
    end
    if (reset) begin // @[GRReg.scala 22:24]
      GRReg_28 <= 64'h0; // @[GRReg.scala 22:24]
    end else if (6'h1c == io_rd_addr[5:0]) begin // @[GRReg.scala 28:23]
      GRReg_28 <= io_ALU_GRReg_IO_rd; // @[GRReg.scala 28:23]
    end
    if (reset) begin // @[GRReg.scala 22:24]
      GRReg_29 <= 64'h0; // @[GRReg.scala 22:24]
    end else if (6'h1d == io_rd_addr[5:0]) begin // @[GRReg.scala 28:23]
      GRReg_29 <= io_ALU_GRReg_IO_rd; // @[GRReg.scala 28:23]
    end
    if (reset) begin // @[GRReg.scala 22:24]
      GRReg_30 <= 64'h0; // @[GRReg.scala 22:24]
    end else if (6'h1e == io_rd_addr[5:0]) begin // @[GRReg.scala 28:23]
      GRReg_30 <= io_ALU_GRReg_IO_rd; // @[GRReg.scala 28:23]
    end
    if (reset) begin // @[GRReg.scala 22:24]
      GRReg_31 <= 64'h0; // @[GRReg.scala 22:24]
    end else if (6'h1f == io_rd_addr[5:0]) begin // @[GRReg.scala 28:23]
      GRReg_31 <= io_ALU_GRReg_IO_rd; // @[GRReg.scala 28:23]
    end
    if (reset) begin // @[GRReg.scala 22:24]
      GRReg_32 <= 64'h0; // @[GRReg.scala 22:24]
    end else if (6'h20 == io_rd_addr[5:0]) begin // @[GRReg.scala 28:23]
      GRReg_32 <= io_ALU_GRReg_IO_rd; // @[GRReg.scala 28:23]
    end
    if (reset) begin // @[GRReg.scala 22:24]
      GRReg_33 <= 64'h0; // @[GRReg.scala 22:24]
    end else if (6'h21 == io_rd_addr[5:0]) begin // @[GRReg.scala 28:23]
      GRReg_33 <= io_ALU_GRReg_IO_rd; // @[GRReg.scala 28:23]
    end
    if (reset) begin // @[GRReg.scala 22:24]
      GRReg_34 <= 64'h0; // @[GRReg.scala 22:24]
    end else if (6'h22 == io_rd_addr[5:0]) begin // @[GRReg.scala 28:23]
      GRReg_34 <= io_ALU_GRReg_IO_rd; // @[GRReg.scala 28:23]
    end
    if (reset) begin // @[GRReg.scala 22:24]
      GRReg_35 <= 64'h0; // @[GRReg.scala 22:24]
    end else if (6'h23 == io_rd_addr[5:0]) begin // @[GRReg.scala 28:23]
      GRReg_35 <= io_ALU_GRReg_IO_rd; // @[GRReg.scala 28:23]
    end
    if (reset) begin // @[GRReg.scala 22:24]
      GRReg_36 <= 64'h0; // @[GRReg.scala 22:24]
    end else if (6'h24 == io_rd_addr[5:0]) begin // @[GRReg.scala 28:23]
      GRReg_36 <= io_ALU_GRReg_IO_rd; // @[GRReg.scala 28:23]
    end
    if (reset) begin // @[GRReg.scala 22:24]
      GRReg_37 <= 64'h0; // @[GRReg.scala 22:24]
    end else if (6'h25 == io_rd_addr[5:0]) begin // @[GRReg.scala 28:23]
      GRReg_37 <= io_ALU_GRReg_IO_rd; // @[GRReg.scala 28:23]
    end
    if (reset) begin // @[GRReg.scala 22:24]
      GRReg_38 <= 64'h0; // @[GRReg.scala 22:24]
    end else if (6'h26 == io_rd_addr[5:0]) begin // @[GRReg.scala 28:23]
      GRReg_38 <= io_ALU_GRReg_IO_rd; // @[GRReg.scala 28:23]
    end
    if (reset) begin // @[GRReg.scala 22:24]
      GRReg_39 <= 64'h0; // @[GRReg.scala 22:24]
    end else if (6'h27 == io_rd_addr[5:0]) begin // @[GRReg.scala 28:23]
      GRReg_39 <= io_ALU_GRReg_IO_rd; // @[GRReg.scala 28:23]
    end
    if (reset) begin // @[GRReg.scala 22:24]
      GRReg_40 <= 64'h0; // @[GRReg.scala 22:24]
    end else if (6'h28 == io_rd_addr[5:0]) begin // @[GRReg.scala 28:23]
      GRReg_40 <= io_ALU_GRReg_IO_rd; // @[GRReg.scala 28:23]
    end
    if (reset) begin // @[GRReg.scala 22:24]
      GRReg_41 <= 64'h0; // @[GRReg.scala 22:24]
    end else if (6'h29 == io_rd_addr[5:0]) begin // @[GRReg.scala 28:23]
      GRReg_41 <= io_ALU_GRReg_IO_rd; // @[GRReg.scala 28:23]
    end
    if (reset) begin // @[GRReg.scala 22:24]
      GRReg_42 <= 64'h0; // @[GRReg.scala 22:24]
    end else if (6'h2a == io_rd_addr[5:0]) begin // @[GRReg.scala 28:23]
      GRReg_42 <= io_ALU_GRReg_IO_rd; // @[GRReg.scala 28:23]
    end
    if (reset) begin // @[GRReg.scala 22:24]
      GRReg_43 <= 64'h0; // @[GRReg.scala 22:24]
    end else if (6'h2b == io_rd_addr[5:0]) begin // @[GRReg.scala 28:23]
      GRReg_43 <= io_ALU_GRReg_IO_rd; // @[GRReg.scala 28:23]
    end
    if (reset) begin // @[GRReg.scala 22:24]
      GRReg_44 <= 64'h0; // @[GRReg.scala 22:24]
    end else if (6'h2c == io_rd_addr[5:0]) begin // @[GRReg.scala 28:23]
      GRReg_44 <= io_ALU_GRReg_IO_rd; // @[GRReg.scala 28:23]
    end
    if (reset) begin // @[GRReg.scala 22:24]
      GRReg_45 <= 64'h0; // @[GRReg.scala 22:24]
    end else if (6'h2d == io_rd_addr[5:0]) begin // @[GRReg.scala 28:23]
      GRReg_45 <= io_ALU_GRReg_IO_rd; // @[GRReg.scala 28:23]
    end
    if (reset) begin // @[GRReg.scala 22:24]
      GRReg_46 <= 64'h0; // @[GRReg.scala 22:24]
    end else if (6'h2e == io_rd_addr[5:0]) begin // @[GRReg.scala 28:23]
      GRReg_46 <= io_ALU_GRReg_IO_rd; // @[GRReg.scala 28:23]
    end
    if (reset) begin // @[GRReg.scala 22:24]
      GRReg_47 <= 64'h0; // @[GRReg.scala 22:24]
    end else if (6'h2f == io_rd_addr[5:0]) begin // @[GRReg.scala 28:23]
      GRReg_47 <= io_ALU_GRReg_IO_rd; // @[GRReg.scala 28:23]
    end
    if (reset) begin // @[GRReg.scala 22:24]
      GRReg_48 <= 64'h0; // @[GRReg.scala 22:24]
    end else if (6'h30 == io_rd_addr[5:0]) begin // @[GRReg.scala 28:23]
      GRReg_48 <= io_ALU_GRReg_IO_rd; // @[GRReg.scala 28:23]
    end
    if (reset) begin // @[GRReg.scala 22:24]
      GRReg_49 <= 64'h0; // @[GRReg.scala 22:24]
    end else if (6'h31 == io_rd_addr[5:0]) begin // @[GRReg.scala 28:23]
      GRReg_49 <= io_ALU_GRReg_IO_rd; // @[GRReg.scala 28:23]
    end
    if (reset) begin // @[GRReg.scala 22:24]
      GRReg_50 <= 64'h0; // @[GRReg.scala 22:24]
    end else if (6'h32 == io_rd_addr[5:0]) begin // @[GRReg.scala 28:23]
      GRReg_50 <= io_ALU_GRReg_IO_rd; // @[GRReg.scala 28:23]
    end
    if (reset) begin // @[GRReg.scala 22:24]
      GRReg_51 <= 64'h0; // @[GRReg.scala 22:24]
    end else if (6'h33 == io_rd_addr[5:0]) begin // @[GRReg.scala 28:23]
      GRReg_51 <= io_ALU_GRReg_IO_rd; // @[GRReg.scala 28:23]
    end
    if (reset) begin // @[GRReg.scala 22:24]
      GRReg_52 <= 64'h0; // @[GRReg.scala 22:24]
    end else if (6'h34 == io_rd_addr[5:0]) begin // @[GRReg.scala 28:23]
      GRReg_52 <= io_ALU_GRReg_IO_rd; // @[GRReg.scala 28:23]
    end
    if (reset) begin // @[GRReg.scala 22:24]
      GRReg_53 <= 64'h0; // @[GRReg.scala 22:24]
    end else if (6'h35 == io_rd_addr[5:0]) begin // @[GRReg.scala 28:23]
      GRReg_53 <= io_ALU_GRReg_IO_rd; // @[GRReg.scala 28:23]
    end
    if (reset) begin // @[GRReg.scala 22:24]
      GRReg_54 <= 64'h0; // @[GRReg.scala 22:24]
    end else if (6'h36 == io_rd_addr[5:0]) begin // @[GRReg.scala 28:23]
      GRReg_54 <= io_ALU_GRReg_IO_rd; // @[GRReg.scala 28:23]
    end
    if (reset) begin // @[GRReg.scala 22:24]
      GRReg_55 <= 64'h0; // @[GRReg.scala 22:24]
    end else if (6'h37 == io_rd_addr[5:0]) begin // @[GRReg.scala 28:23]
      GRReg_55 <= io_ALU_GRReg_IO_rd; // @[GRReg.scala 28:23]
    end
    if (reset) begin // @[GRReg.scala 22:24]
      GRReg_56 <= 64'h0; // @[GRReg.scala 22:24]
    end else if (6'h38 == io_rd_addr[5:0]) begin // @[GRReg.scala 28:23]
      GRReg_56 <= io_ALU_GRReg_IO_rd; // @[GRReg.scala 28:23]
    end
    if (reset) begin // @[GRReg.scala 22:24]
      GRReg_57 <= 64'h0; // @[GRReg.scala 22:24]
    end else if (6'h39 == io_rd_addr[5:0]) begin // @[GRReg.scala 28:23]
      GRReg_57 <= io_ALU_GRReg_IO_rd; // @[GRReg.scala 28:23]
    end
    if (reset) begin // @[GRReg.scala 22:24]
      GRReg_58 <= 64'h0; // @[GRReg.scala 22:24]
    end else if (6'h3a == io_rd_addr[5:0]) begin // @[GRReg.scala 28:23]
      GRReg_58 <= io_ALU_GRReg_IO_rd; // @[GRReg.scala 28:23]
    end
    if (reset) begin // @[GRReg.scala 22:24]
      GRReg_59 <= 64'h0; // @[GRReg.scala 22:24]
    end else if (6'h3b == io_rd_addr[5:0]) begin // @[GRReg.scala 28:23]
      GRReg_59 <= io_ALU_GRReg_IO_rd; // @[GRReg.scala 28:23]
    end
    if (reset) begin // @[GRReg.scala 22:24]
      GRReg_60 <= 64'h0; // @[GRReg.scala 22:24]
    end else if (6'h3c == io_rd_addr[5:0]) begin // @[GRReg.scala 28:23]
      GRReg_60 <= io_ALU_GRReg_IO_rd; // @[GRReg.scala 28:23]
    end
    if (reset) begin // @[GRReg.scala 22:24]
      GRReg_61 <= 64'h0; // @[GRReg.scala 22:24]
    end else if (6'h3d == io_rd_addr[5:0]) begin // @[GRReg.scala 28:23]
      GRReg_61 <= io_ALU_GRReg_IO_rd; // @[GRReg.scala 28:23]
    end
    if (reset) begin // @[GRReg.scala 22:24]
      GRReg_62 <= 64'h0; // @[GRReg.scala 22:24]
    end else if (6'h3e == io_rd_addr[5:0]) begin // @[GRReg.scala 28:23]
      GRReg_62 <= io_ALU_GRReg_IO_rd; // @[GRReg.scala 28:23]
    end
    if (reset) begin // @[GRReg.scala 22:24]
      GRReg_63 <= 64'h0; // @[GRReg.scala 22:24]
    end else if (6'h3f == io_rd_addr[5:0]) begin // @[GRReg.scala 28:23]
      GRReg_63 <= io_ALU_GRReg_IO_rd; // @[GRReg.scala 28:23]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  GRReg_0 = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  GRReg_1 = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  GRReg_2 = _RAND_2[63:0];
  _RAND_3 = {2{`RANDOM}};
  GRReg_3 = _RAND_3[63:0];
  _RAND_4 = {2{`RANDOM}};
  GRReg_4 = _RAND_4[63:0];
  _RAND_5 = {2{`RANDOM}};
  GRReg_5 = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  GRReg_6 = _RAND_6[63:0];
  _RAND_7 = {2{`RANDOM}};
  GRReg_7 = _RAND_7[63:0];
  _RAND_8 = {2{`RANDOM}};
  GRReg_8 = _RAND_8[63:0];
  _RAND_9 = {2{`RANDOM}};
  GRReg_9 = _RAND_9[63:0];
  _RAND_10 = {2{`RANDOM}};
  GRReg_10 = _RAND_10[63:0];
  _RAND_11 = {2{`RANDOM}};
  GRReg_11 = _RAND_11[63:0];
  _RAND_12 = {2{`RANDOM}};
  GRReg_12 = _RAND_12[63:0];
  _RAND_13 = {2{`RANDOM}};
  GRReg_13 = _RAND_13[63:0];
  _RAND_14 = {2{`RANDOM}};
  GRReg_14 = _RAND_14[63:0];
  _RAND_15 = {2{`RANDOM}};
  GRReg_15 = _RAND_15[63:0];
  _RAND_16 = {2{`RANDOM}};
  GRReg_16 = _RAND_16[63:0];
  _RAND_17 = {2{`RANDOM}};
  GRReg_17 = _RAND_17[63:0];
  _RAND_18 = {2{`RANDOM}};
  GRReg_18 = _RAND_18[63:0];
  _RAND_19 = {2{`RANDOM}};
  GRReg_19 = _RAND_19[63:0];
  _RAND_20 = {2{`RANDOM}};
  GRReg_20 = _RAND_20[63:0];
  _RAND_21 = {2{`RANDOM}};
  GRReg_21 = _RAND_21[63:0];
  _RAND_22 = {2{`RANDOM}};
  GRReg_22 = _RAND_22[63:0];
  _RAND_23 = {2{`RANDOM}};
  GRReg_23 = _RAND_23[63:0];
  _RAND_24 = {2{`RANDOM}};
  GRReg_24 = _RAND_24[63:0];
  _RAND_25 = {2{`RANDOM}};
  GRReg_25 = _RAND_25[63:0];
  _RAND_26 = {2{`RANDOM}};
  GRReg_26 = _RAND_26[63:0];
  _RAND_27 = {2{`RANDOM}};
  GRReg_27 = _RAND_27[63:0];
  _RAND_28 = {2{`RANDOM}};
  GRReg_28 = _RAND_28[63:0];
  _RAND_29 = {2{`RANDOM}};
  GRReg_29 = _RAND_29[63:0];
  _RAND_30 = {2{`RANDOM}};
  GRReg_30 = _RAND_30[63:0];
  _RAND_31 = {2{`RANDOM}};
  GRReg_31 = _RAND_31[63:0];
  _RAND_32 = {2{`RANDOM}};
  GRReg_32 = _RAND_32[63:0];
  _RAND_33 = {2{`RANDOM}};
  GRReg_33 = _RAND_33[63:0];
  _RAND_34 = {2{`RANDOM}};
  GRReg_34 = _RAND_34[63:0];
  _RAND_35 = {2{`RANDOM}};
  GRReg_35 = _RAND_35[63:0];
  _RAND_36 = {2{`RANDOM}};
  GRReg_36 = _RAND_36[63:0];
  _RAND_37 = {2{`RANDOM}};
  GRReg_37 = _RAND_37[63:0];
  _RAND_38 = {2{`RANDOM}};
  GRReg_38 = _RAND_38[63:0];
  _RAND_39 = {2{`RANDOM}};
  GRReg_39 = _RAND_39[63:0];
  _RAND_40 = {2{`RANDOM}};
  GRReg_40 = _RAND_40[63:0];
  _RAND_41 = {2{`RANDOM}};
  GRReg_41 = _RAND_41[63:0];
  _RAND_42 = {2{`RANDOM}};
  GRReg_42 = _RAND_42[63:0];
  _RAND_43 = {2{`RANDOM}};
  GRReg_43 = _RAND_43[63:0];
  _RAND_44 = {2{`RANDOM}};
  GRReg_44 = _RAND_44[63:0];
  _RAND_45 = {2{`RANDOM}};
  GRReg_45 = _RAND_45[63:0];
  _RAND_46 = {2{`RANDOM}};
  GRReg_46 = _RAND_46[63:0];
  _RAND_47 = {2{`RANDOM}};
  GRReg_47 = _RAND_47[63:0];
  _RAND_48 = {2{`RANDOM}};
  GRReg_48 = _RAND_48[63:0];
  _RAND_49 = {2{`RANDOM}};
  GRReg_49 = _RAND_49[63:0];
  _RAND_50 = {2{`RANDOM}};
  GRReg_50 = _RAND_50[63:0];
  _RAND_51 = {2{`RANDOM}};
  GRReg_51 = _RAND_51[63:0];
  _RAND_52 = {2{`RANDOM}};
  GRReg_52 = _RAND_52[63:0];
  _RAND_53 = {2{`RANDOM}};
  GRReg_53 = _RAND_53[63:0];
  _RAND_54 = {2{`RANDOM}};
  GRReg_54 = _RAND_54[63:0];
  _RAND_55 = {2{`RANDOM}};
  GRReg_55 = _RAND_55[63:0];
  _RAND_56 = {2{`RANDOM}};
  GRReg_56 = _RAND_56[63:0];
  _RAND_57 = {2{`RANDOM}};
  GRReg_57 = _RAND_57[63:0];
  _RAND_58 = {2{`RANDOM}};
  GRReg_58 = _RAND_58[63:0];
  _RAND_59 = {2{`RANDOM}};
  GRReg_59 = _RAND_59[63:0];
  _RAND_60 = {2{`RANDOM}};
  GRReg_60 = _RAND_60[63:0];
  _RAND_61 = {2{`RANDOM}};
  GRReg_61 = _RAND_61[63:0];
  _RAND_62 = {2{`RANDOM}};
  GRReg_62 = _RAND_62[63:0];
  _RAND_63 = {2{`RANDOM}};
  GRReg_63 = _RAND_63[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
