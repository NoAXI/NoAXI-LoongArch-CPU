module ALU(
  input         clock,
  input         reset,
  input  [31:0] io_instruction,
  input  [63:0] io_rj,
  input  [63:0] io_rk,
  input  [63:0] io_rd_in,
  input  [63:0] io_imm,
  output [63:0] io_rd
);
  wire [31:0] _T = io_instruction & 32'h1ffff000; // @[ALU.scala 27:26]
  wire [31:0] _io_rd_T_3 = io_rj[31:0] + io_rk[31:0]; // @[ALU.scala 28:44]
  wire [31:0] io_rd_fill = _io_rd_T_3[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 74:12]
  wire [63:0] _io_rd_T_4 = {io_rd_fill,_io_rd_T_3}; // @[Cat.scala 31:58]
  wire [63:0] _io_rd_T_6 = io_rj + io_rk; // @[ALU.scala 30:24]
  wire [31:0] _io_rd_T_10 = io_rj[31:0] - io_rk[31:0]; // @[ALU.scala 32:44]
  wire [31:0] io_rd_fill_1 = _io_rd_T_10[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 74:12]
  wire [63:0] _io_rd_T_11 = {io_rd_fill_1,_io_rd_T_10}; // @[Cat.scala 31:58]
  wire [63:0] _io_rd_T_13 = io_rj - io_rk; // @[ALU.scala 34:24]
  wire [31:0] _T_8 = io_instruction & 32'h1ff80000; // @[ALU.scala 35:33]
  wire [19:0] io_rd_fill_2 = io_imm[11] ? 20'hfffff : 20'h0; // @[Bitwise.scala 74:12]
  wire [31:0] _io_rd_T_16 = {io_rd_fill_2,io_imm[11:0]}; // @[Cat.scala 31:58]
  wire [31:0] _io_rd_T_18 = io_rj[31:0] + _io_rd_T_16; // @[ALU.scala 36:44]
  wire [31:0] io_rd_fill_3 = _io_rd_T_18[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 74:12]
  wire [63:0] _io_rd_T_19 = {io_rd_fill_3,_io_rd_T_18}; // @[Cat.scala 31:58]
  wire [51:0] io_rd_fill_4 = io_imm[11] ? 52'hfffffffffffff : 52'h0; // @[Bitwise.scala 74:12]
  wire [63:0] _io_rd_T_21 = {io_rd_fill_4,io_imm[11:0]}; // @[Cat.scala 31:58]
  wire [63:0] _io_rd_T_23 = io_rj + _io_rd_T_21; // @[ALU.scala 39:24]
  wire [31:0] _T_12 = io_instruction & 32'h1f800000; // @[ALU.scala 40:33]
  wire [31:0] _io_rd_T_26 = {io_imm[15:0],16'h0}; // @[Cat.scala 31:58]
  wire [31:0] io_rd_fill_5 = _io_rd_T_26[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 74:12]
  wire [63:0] _io_rd_T_27 = {io_rd_fill_5,io_imm[15:0],16'h0}; // @[Cat.scala 31:58]
  wire [63:0] _io_rd_T_29 = io_rj + _io_rd_T_27; // @[ALU.scala 41:24]
  wire [31:0] _T_14 = io_instruction & 32'h1fffc000; // @[ALU.scala 42:33]
  wire [1:0] _io_rd_T_33 = io_imm[1:0] + 2'h1; // @[ALU.scala 43:62]
  wire [34:0] _GEN_14 = {{3'd0}, io_rj[31:0]}; // @[ALU.scala 43:45]
  wire [34:0] _io_rd_T_34 = _GEN_14 << _io_rd_T_33; // @[ALU.scala 43:45]
  wire [34:0] _GEN_13 = {{3'd0}, io_rk[31:0]}; // @[ALU.scala 43:70]
  wire [34:0] _io_rd_T_37 = _io_rd_T_34 + _GEN_13; // @[ALU.scala 43:70]
  wire [28:0] io_rd_fill_6 = _io_rd_T_37[34] ? 29'h1fffffff : 29'h0; // @[Bitwise.scala 74:12]
  wire [63:0] _io_rd_T_38 = {io_rd_fill_6,_io_rd_T_37}; // @[Cat.scala 31:58]
  wire [63:0] _io_rd_T_47 = {29'h0,_io_rd_T_37}; // @[Cat.scala 31:58]
  wire [31:0] _T_18 = io_instruction & 32'h1fff8000; // @[ALU.scala 46:33]
  wire [66:0] _GEN_16 = {{3'd0}, io_rj}; // @[ALU.scala 47:25]
  wire [66:0] _io_rd_T_51 = _GEN_16 << _io_rd_T_33; // @[ALU.scala 47:25]
  wire [66:0] _GEN_15 = {{3'd0}, io_rk}; // @[ALU.scala 47:50]
  wire [66:0] _io_rd_T_53 = _io_rd_T_51 + _GEN_15; // @[ALU.scala 47:50]
  wire [31:0] _T_20 = io_instruction & 32'h1fc00000; // @[ALU.scala 48:33]
  wire [31:0] _io_rd_T_56 = {io_imm[19:0],12'h0}; // @[Cat.scala 31:58]
  wire [31:0] io_rd_fill_8 = _io_rd_T_56[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 74:12]
  wire [63:0] _io_rd_T_57 = {io_rd_fill_8,io_imm[19:0],12'h0}; // @[Cat.scala 31:58]
  wire [11:0] io_rd_fill_9 = io_imm[19] ? 12'hfff : 12'h0; // @[Bitwise.scala 74:12]
  wire [63:0] _io_rd_T_61 = {io_rd_fill_9,io_imm[19:0],io_rd_in[31:0]}; // @[Cat.scala 31:58]
  wire [63:0] _io_rd_T_64 = {io_imm[11:0],io_rj[51:0]}; // @[Cat.scala 31:58]
  wire [63:0] _GEN_0 = 32'h600000 == _T_8 ? _io_rd_T_64 : 64'h0; // @[ALU.scala 25:11 52:46 53:15]
  wire [63:0] _GEN_1 = 32'h2c00000 == _T_20 ? _io_rd_T_61 : _GEN_0; // @[ALU.scala 50:46 51:15]
  wire [63:0] _GEN_2 = 32'h2800000 == _T_20 ? _io_rd_T_57 : _GEN_1; // @[ALU.scala 48:46 49:15]
  wire [66:0] _GEN_3 = 32'h58000 == _T_18 ? _io_rd_T_53 : {{3'd0}, _GEN_2}; // @[ALU.scala 46:45 47:15]
  wire [66:0] _GEN_4 = 32'hc000 == _T_14 ? {{3'd0}, _io_rd_T_47} : _GEN_3; // @[ALU.scala 44:46 45:15]
  wire [66:0] _GEN_5 = 32'h8000 == _T_14 ? {{3'd0}, _io_rd_T_38} : _GEN_4; // @[ALU.scala 42:45 43:15]
  wire [66:0] _GEN_6 = 32'h2000000 == _T_12 ? {{3'd0}, _io_rd_T_29} : _GEN_5; // @[ALU.scala 40:48 41:15]
  wire [66:0] _GEN_7 = 32'h580000 == _T_8 ? {{3'd0}, _io_rd_T_23} : _GEN_6; // @[ALU.scala 38:45 39:15]
  wire [66:0] _GEN_8 = 32'h500000 == _T_8 ? {{3'd0}, _io_rd_T_19} : _GEN_7; // @[ALU.scala 35:45 36:15]
  wire [66:0] _GEN_9 = 32'h23000 == _T ? {{3'd0}, _io_rd_T_13} : _GEN_8; // @[ALU.scala 33:44 34:15]
  wire [66:0] _GEN_10 = 32'h22000 == _T ? {{3'd0}, _io_rd_T_11} : _GEN_9; // @[ALU.scala 31:44 32:15]
  wire [66:0] _GEN_11 = 32'h21000 == _T ? {{3'd0}, _io_rd_T_6} : _GEN_10; // @[ALU.scala 29:44 30:15]
  wire [66:0] _GEN_12 = 32'h20000 == _T ? {{3'd0}, _io_rd_T_4} : _GEN_11; // @[ALU.scala 27:37 28:15]
  assign io_rd = _GEN_12[63:0];
endmodule
